I-D vs V_DS

.include ALD1105P.txt

m1 1 2 0 0 ALD1105P
vgg 3 0 dc -5V
r2 4 0 1.5k
r1 3 4 3.5k
r3 3 5 4.7k
r4 5 0 200
vdummy1 1 5 dc 0V
vdummy2 2 4 dc 0V 

.dc r2 1 5k 0.1

.control
run

plot i(vdummy1) vs v(2)

set hcopydevtype = postscript
set hcopypscolor = 1
hardcopy Part1_P i(vdummy1) vs v(2)

.endc
.end
